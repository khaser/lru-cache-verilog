module cache(clk, c_dump, reset);


endmodule
