module cpu(out, in1, in2);


endmodule
